
module current_state ( ph1, ph2, regwrite, reset, ra, wa, wd, rd );
  input [2:0] ra;
  input [2:0] wa;
  input [7:0] wd;
  output [7:0] rd;
  input ph1, ph2, regwrite, reset;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, N27, N28, N31, N36, N37, N38,
         N39, N40, N41, N42, N43, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77;
  wire   [63:0] RAM;

  latch_c_1x RAM_reg_7__7_ ( .ph(N43), .d(N25), .q(RAM[63]) );
  latch_c_1x RAM_reg_7__6_ ( .ph(N43), .d(N24), .q(RAM[62]) );
  latch_c_1x RAM_reg_7__5_ ( .ph(N43), .d(N23), .q(RAM[61]) );
  latch_c_1x RAM_reg_7__4_ ( .ph(N43), .d(N31), .q(RAM[60]) );
  latch_c_1x RAM_reg_7__3_ ( .ph(N43), .d(N27), .q(RAM[59]) );
  latch_c_1x RAM_reg_7__2_ ( .ph(N43), .d(N20), .q(RAM[58]) );
  latch_c_1x RAM_reg_7__1_ ( .ph(N43), .d(N19), .q(RAM[57]) );
  latch_c_1x RAM_reg_7__0_ ( .ph(N43), .d(N18), .q(RAM[56]) );
  latch_c_1x RAM_reg_6__7_ ( .ph(N42), .d(N25), .q(RAM[55]) );
  latch_c_1x RAM_reg_6__6_ ( .ph(N42), .d(N24), .q(RAM[54]) );
  latch_c_1x RAM_reg_6__5_ ( .ph(N42), .d(N23), .q(RAM[53]) );
  latch_c_1x RAM_reg_6__4_ ( .ph(N42), .d(N31), .q(RAM[52]) );
  latch_c_1x RAM_reg_6__3_ ( .ph(N42), .d(N27), .q(RAM[51]) );
  latch_c_1x RAM_reg_6__2_ ( .ph(N42), .d(N20), .q(RAM[50]) );
  latch_c_1x RAM_reg_6__1_ ( .ph(N42), .d(N19), .q(RAM[49]) );
  latch_c_1x RAM_reg_6__0_ ( .ph(N42), .d(N18), .q(RAM[48]) );
  latch_c_1x RAM_reg_5__7_ ( .ph(N41), .d(N25), .q(RAM[47]) );
  latch_c_1x RAM_reg_5__6_ ( .ph(N41), .d(N24), .q(RAM[46]) );
  latch_c_1x RAM_reg_5__5_ ( .ph(N41), .d(N23), .q(RAM[45]) );
  latch_c_1x RAM_reg_5__4_ ( .ph(N41), .d(N31), .q(RAM[44]) );
  latch_c_1x RAM_reg_5__3_ ( .ph(N41), .d(N27), .q(RAM[43]) );
  latch_c_1x RAM_reg_5__2_ ( .ph(N41), .d(N20), .q(RAM[42]) );
  latch_c_1x RAM_reg_5__1_ ( .ph(N41), .d(N19), .q(RAM[41]) );
  latch_c_1x RAM_reg_5__0_ ( .ph(N41), .d(N18), .q(RAM[40]) );
  latch_c_1x RAM_reg_4__7_ ( .ph(N40), .d(N25), .q(RAM[39]) );
  latch_c_1x RAM_reg_4__6_ ( .ph(N40), .d(N24), .q(RAM[38]) );
  latch_c_1x RAM_reg_4__5_ ( .ph(N40), .d(N23), .q(RAM[37]) );
  latch_c_1x RAM_reg_4__4_ ( .ph(N40), .d(N31), .q(RAM[36]) );
  latch_c_1x RAM_reg_4__3_ ( .ph(N40), .d(N27), .q(RAM[35]) );
  latch_c_1x RAM_reg_4__2_ ( .ph(N40), .d(N20), .q(RAM[34]) );
  latch_c_1x RAM_reg_4__1_ ( .ph(N40), .d(N19), .q(RAM[33]) );
  latch_c_1x RAM_reg_4__0_ ( .ph(N40), .d(N18), .q(RAM[32]) );
  latch_c_1x RAM_reg_3__7_ ( .ph(N39), .d(N25), .q(RAM[31]) );
  latch_c_1x RAM_reg_3__6_ ( .ph(N39), .d(N24), .q(RAM[30]) );
  latch_c_1x RAM_reg_3__5_ ( .ph(N39), .d(N23), .q(RAM[29]) );
  latch_c_1x RAM_reg_3__4_ ( .ph(N39), .d(N31), .q(RAM[28]) );
  latch_c_1x RAM_reg_3__3_ ( .ph(N39), .d(N27), .q(RAM[27]) );
  latch_c_1x RAM_reg_3__2_ ( .ph(N39), .d(N20), .q(RAM[26]) );
  latch_c_1x RAM_reg_3__1_ ( .ph(N39), .d(N19), .q(RAM[25]) );
  latch_c_1x RAM_reg_3__0_ ( .ph(N39), .d(N18), .q(RAM[24]) );
  latch_c_1x RAM_reg_2__7_ ( .ph(N38), .d(N25), .q(RAM[23]) );
  latch_c_1x RAM_reg_2__6_ ( .ph(N38), .d(N24), .q(RAM[22]) );
  latch_c_1x RAM_reg_2__5_ ( .ph(N38), .d(N23), .q(RAM[21]) );
  latch_c_1x RAM_reg_2__4_ ( .ph(N38), .d(N22), .q(RAM[20]) );
  latch_c_1x RAM_reg_2__3_ ( .ph(N38), .d(N27), .q(RAM[19]) );
  latch_c_1x RAM_reg_2__2_ ( .ph(N38), .d(N20), .q(RAM[18]) );
  latch_c_1x RAM_reg_2__1_ ( .ph(N38), .d(N19), .q(RAM[17]) );
  latch_c_1x RAM_reg_2__0_ ( .ph(N38), .d(N18), .q(RAM[16]) );
  latch_c_1x RAM_reg_1__7_ ( .ph(N37), .d(N25), .q(RAM[15]) );
  latch_c_1x RAM_reg_1__6_ ( .ph(N37), .d(N24), .q(RAM[14]) );
  latch_c_1x RAM_reg_1__5_ ( .ph(N37), .d(N28), .q(RAM[13]) );
  latch_c_1x RAM_reg_1__4_ ( .ph(N37), .d(N22), .q(RAM[12]) );
  latch_c_1x RAM_reg_1__3_ ( .ph(N37), .d(N27), .q(RAM[11]) );
  latch_c_1x RAM_reg_1__2_ ( .ph(N37), .d(N20), .q(RAM[10]) );
  latch_c_1x RAM_reg_1__1_ ( .ph(N37), .d(N19), .q(RAM[9]) );
  latch_c_1x RAM_reg_1__0_ ( .ph(N37), .d(N18), .q(RAM[8]) );
  latch_c_1x RAM_reg_0__7_ ( .ph(N36), .d(N25), .q(RAM[7]) );
  latch_c_1x RAM_reg_0__6_ ( .ph(N36), .d(N24), .q(RAM[6]) );
  latch_c_1x RAM_reg_0__5_ ( .ph(N36), .d(N23), .q(RAM[5]) );
  latch_c_1x RAM_reg_0__4_ ( .ph(N36), .d(N22), .q(RAM[4]) );
  latch_c_1x RAM_reg_0__3_ ( .ph(N36), .d(N21), .q(RAM[3]) );
  latch_c_1x RAM_reg_0__2_ ( .ph(N36), .d(N20), .q(RAM[2]) );
  latch_c_1x RAM_reg_0__1_ ( .ph(N36), .d(N19), .q(RAM[1]) );
  latch_c_1x RAM_reg_0__0_ ( .ph(N36), .d(N18), .q(RAM[0]) );
  inv_4x U35 ( .a(reset), .y(n17) );
  nor2_1x U36 ( .a(n23), .b(n22), .y(n28) );
  nor2_1x U37 ( .a(wa[2]), .b(n22), .y(n21) );
  nand2_1x U38 ( .a(ph2), .b(n18), .y(n22) );
  nor2_1x U39 ( .a(n20), .b(n19), .y(n29) );
  nor2_1x U40 ( .a(wa[1]), .b(n19), .y(n25) );
  inv_1x U41 ( .a(wa[0]), .y(n19) );
  inv_1x U42 ( .a(wa[1]), .y(n20) );
  inv_1x U43 ( .a(wa[2]), .y(n23) );
  nor2_2x U44 ( .a(wa[0]), .b(n20), .y(n26) );
  nor2_2x U45 ( .a(wa[1]), .b(wa[0]), .y(n24) );
  inv_4x U46 ( .a(n15), .y(N31) );
  nand2_2x U47 ( .a(n17), .b(n16), .y(N28) );
  inv_4x U48 ( .a(n14), .y(N27) );
  nand2_2x U49 ( .a(n17), .b(n14), .y(N21) );
  nand2_1x U50 ( .a(n18), .b(wd[3]), .y(n14) );
  inv_4x U51 ( .a(n16), .y(N23) );
  nand2_1x U52 ( .a(n18), .b(wd[5]), .y(n16) );
  nand2_2x U53 ( .a(n17), .b(n15), .y(N22) );
  and2_1x U54 ( .a(regwrite), .b(n17), .y(n18) );
  and2_1x U55 ( .a(n18), .b(wd[0]), .y(N18) );
  and2_1x U56 ( .a(n18), .b(wd[1]), .y(N19) );
  and2_1x U57 ( .a(n18), .b(wd[2]), .y(N20) );
  nand2_1x U58 ( .a(n18), .b(wd[4]), .y(n15) );
  and2_1x U59 ( .a(n18), .b(wd[6]), .y(N24) );
  and2_1x U60 ( .a(n18), .b(wd[7]), .y(N25) );
  and2_1x U61 ( .a(reset), .b(ph2), .y(n27) );
  a2o1_1x U62 ( .a(n24), .b(n21), .c(n27), .y(N36) );
  a2o1_1x U63 ( .a(n21), .b(n25), .c(n27), .y(N37) );
  a2o1_1x U64 ( .a(n21), .b(n26), .c(n27), .y(N38) );
  a2o1_1x U65 ( .a(n21), .b(n29), .c(n27), .y(N39) );
  a2o1_1x U66 ( .a(n24), .b(n28), .c(n27), .y(N40) );
  a2o1_1x U67 ( .a(n25), .b(n28), .c(n27), .y(N41) );
  a2o1_1x U68 ( .a(n26), .b(n28), .c(n27), .y(N42) );
  a2o1_1x U69 ( .a(n29), .b(n28), .c(n27), .y(N43) );
  mux2_c_1x U70 ( .d0(RAM[0]), .d1(RAM[8]), .s(ra[0]), .y(n30) );
  mux2_c_1x U71 ( .d0(RAM[16]), .d1(RAM[24]), .s(ra[0]), .y(n31) );
  mux2_c_1x U72 ( .d0(RAM[32]), .d1(RAM[40]), .s(ra[0]), .y(n32) );
  mux2_c_1x U73 ( .d0(RAM[48]), .d1(RAM[56]), .s(ra[0]), .y(n33) );
  mux2_c_1x U74 ( .d0(n30), .d1(n31), .s(ra[1]), .y(n34) );
  mux2_c_1x U75 ( .d0(n32), .d1(n33), .s(ra[1]), .y(n35) );
  mux2_c_1x U76 ( .d0(n34), .d1(n35), .s(ra[2]), .y(rd[0]) );
  mux2_c_1x U77 ( .d0(RAM[1]), .d1(RAM[9]), .s(ra[0]), .y(n36) );
  mux2_c_1x U78 ( .d0(RAM[17]), .d1(RAM[25]), .s(ra[0]), .y(n37) );
  mux2_c_1x U79 ( .d0(RAM[33]), .d1(RAM[41]), .s(ra[0]), .y(n38) );
  mux2_c_1x U80 ( .d0(RAM[49]), .d1(RAM[57]), .s(ra[0]), .y(n39) );
  mux2_c_1x U81 ( .d0(n36), .d1(n37), .s(ra[1]), .y(n40) );
  mux2_c_1x U82 ( .d0(n38), .d1(n39), .s(ra[1]), .y(n41) );
  mux2_c_1x U83 ( .d0(n40), .d1(n41), .s(ra[2]), .y(rd[1]) );
  mux2_c_1x U84 ( .d0(RAM[2]), .d1(RAM[10]), .s(ra[0]), .y(n42) );
  mux2_c_1x U85 ( .d0(RAM[18]), .d1(RAM[26]), .s(ra[0]), .y(n43) );
  mux2_c_1x U86 ( .d0(RAM[34]), .d1(RAM[42]), .s(ra[0]), .y(n44) );
  mux2_c_1x U87 ( .d0(RAM[50]), .d1(RAM[58]), .s(ra[0]), .y(n45) );
  mux2_c_1x U88 ( .d0(n42), .d1(n43), .s(ra[1]), .y(n46) );
  mux2_c_1x U89 ( .d0(n44), .d1(n45), .s(ra[1]), .y(n47) );
  mux2_c_1x U90 ( .d0(n46), .d1(n47), .s(ra[2]), .y(rd[2]) );
  mux2_c_1x U91 ( .d0(RAM[3]), .d1(RAM[11]), .s(ra[0]), .y(n48) );
  mux2_c_1x U92 ( .d0(RAM[19]), .d1(RAM[27]), .s(ra[0]), .y(n49) );
  mux2_c_1x U93 ( .d0(RAM[35]), .d1(RAM[43]), .s(ra[0]), .y(n50) );
  mux2_c_1x U94 ( .d0(RAM[51]), .d1(RAM[59]), .s(ra[0]), .y(n51) );
  mux2_c_1x U95 ( .d0(n48), .d1(n49), .s(ra[1]), .y(n52) );
  mux2_c_1x U96 ( .d0(n50), .d1(n51), .s(ra[1]), .y(n53) );
  mux2_c_1x U97 ( .d0(n52), .d1(n53), .s(ra[2]), .y(rd[3]) );
  mux2_c_1x U98 ( .d0(RAM[4]), .d1(RAM[12]), .s(ra[0]), .y(n54) );
  mux2_c_1x U99 ( .d0(RAM[20]), .d1(RAM[28]), .s(ra[0]), .y(n55) );
  mux2_c_1x U100 ( .d0(RAM[36]), .d1(RAM[44]), .s(ra[0]), .y(n56) );
  mux2_c_1x U101 ( .d0(RAM[52]), .d1(RAM[60]), .s(ra[0]), .y(n57) );
  mux2_c_1x U102 ( .d0(n54), .d1(n55), .s(ra[1]), .y(n58) );
  mux2_c_1x U103 ( .d0(n56), .d1(n57), .s(ra[1]), .y(n59) );
  mux2_c_1x U104 ( .d0(n58), .d1(n59), .s(ra[2]), .y(rd[4]) );
  mux2_c_1x U105 ( .d0(RAM[5]), .d1(RAM[13]), .s(ra[0]), .y(n60) );
  mux2_c_1x U106 ( .d0(RAM[21]), .d1(RAM[29]), .s(ra[0]), .y(n61) );
  mux2_c_1x U107 ( .d0(RAM[37]), .d1(RAM[45]), .s(ra[0]), .y(n62) );
  mux2_c_1x U108 ( .d0(RAM[53]), .d1(RAM[61]), .s(ra[0]), .y(n63) );
  mux2_c_1x U109 ( .d0(n60), .d1(n61), .s(ra[1]), .y(n64) );
  mux2_c_1x U110 ( .d0(n62), .d1(n63), .s(ra[1]), .y(n65) );
  mux2_c_1x U111 ( .d0(n64), .d1(n65), .s(ra[2]), .y(rd[5]) );
  mux2_c_1x U112 ( .d0(RAM[6]), .d1(RAM[14]), .s(ra[0]), .y(n66) );
  mux2_c_1x U113 ( .d0(RAM[22]), .d1(RAM[30]), .s(ra[0]), .y(n67) );
  mux2_c_1x U114 ( .d0(RAM[38]), .d1(RAM[46]), .s(ra[0]), .y(n68) );
  mux2_c_1x U115 ( .d0(RAM[54]), .d1(RAM[62]), .s(ra[0]), .y(n69) );
  mux2_c_1x U116 ( .d0(n66), .d1(n67), .s(ra[1]), .y(n70) );
  mux2_c_1x U117 ( .d0(n68), .d1(n69), .s(ra[1]), .y(n71) );
  mux2_c_1x U118 ( .d0(n70), .d1(n71), .s(ra[2]), .y(rd[6]) );
  mux2_c_1x U119 ( .d0(RAM[7]), .d1(RAM[15]), .s(ra[0]), .y(n72) );
  mux2_c_1x U120 ( .d0(RAM[23]), .d1(RAM[31]), .s(ra[0]), .y(n73) );
  mux2_c_1x U121 ( .d0(RAM[39]), .d1(RAM[47]), .s(ra[0]), .y(n74) );
  mux2_c_1x U122 ( .d0(RAM[55]), .d1(RAM[63]), .s(ra[0]), .y(n75) );
  mux2_c_1x U123 ( .d0(n72), .d1(n73), .s(ra[1]), .y(n76) );
  mux2_c_1x U124 ( .d0(n74), .d1(n75), .s(ra[1]), .y(n77) );
  mux2_c_1x U125 ( .d0(n76), .d1(n77), .s(ra[2]), .y(rd[7]) );
endmodule

